module Dispatch (

);

endmodule
