module Issue (

);

endmodule
