module VTop (

);

endmodule
