module Adder (

);

endmodule
