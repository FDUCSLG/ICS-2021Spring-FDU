`ifndef __OOO_DEFS_SVH__
`define __OOO_DEFS_SVH__

// verilator lint_save
// verilator lint_off UNUSED

parameter int N_ISSUE_ENTRIES    = 4;
parameter int N_DISPATCH_ENTRIES = 2;
parameter int N_COMMIT_ENTRIES   = 8;

// verilator lint_restore

`endif
