module Mult (

);

endmodule
