module RegisterFile (

);

endmodule
